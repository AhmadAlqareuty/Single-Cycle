module ahmad();
endmodule